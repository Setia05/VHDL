library IEEE;
use IEEE.std_logic_1164.all;
 
entity nor_gate is
Port( A : in std_logic;
		B : in std_logic;
		C : in std_logic;
		Y : out std_logic);
end nor_gate;
architecture Behavioral of and_gate is
begin

	Y<=(A nor B);
	
end Behavioral;
